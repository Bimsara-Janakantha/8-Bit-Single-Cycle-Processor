/*
    * CO224 - Computer Architecture
    * Lab 05 - Part 5
    * and unit
    * Group 09 (E/20/148, E/20/157)
    * 2024-05-15
    * Version 1.0
*/

`timescale 1ns/100ps

// ALU and unit is used to do and operation in the ALU
module myAND(DATA1, DATA2, RESULT);
    // Input-output Declaration
    input [7:0] DATA1, DATA2;
    output [7:0] RESULT;

    // Result
    assign #1 RESULT = DATA1 & DATA2;
endmodule